// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package ibex_rvfi_pkg;
  import uvm_pkg::*;

  `include "uvm_macros.svh"

  `include "ibex_rvfi_seq_item.sv"
  `include "ibex_rvfi_monitor.sv"
endpackage
