package core_ibex_testrig_env_pkg;
  import uvm_pkg::*;
  import ibex_testrig_agent_pkg::*;

  `include "uvm_macros.svh"

  `include "core_ibex_testrig_env.sv"
endpackage
