// Copyright lowRISC contributors.
// Licensed under the Apache License, Version 2.0, see LICENSE for details.
// SPDX-License-Identifier: Apache-2.0

package ibex_testrig_agent_pkg;
  import uvm_pkg::*;
  import ibex_rvfi_pkg::*;

  `include "uvm_macros.svh"

  `include "testrig_dpi.svh"
  `include "ibex_testrig_dii_driver.sv"
  `include "ibex_testrig_agent.sv"
endpackage
